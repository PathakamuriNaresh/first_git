this is the file created in the sub1 branch
this is the first time modified
