this is the file created in the sub1 branch
